`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08/03/2021 08:46:43 PM
// Design Name: 
// Module Name: Miner
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

/*
TODO:
	Replace integers for reg
	Combine hashValues and oldHashValues into array
	Create target check
	Improve Choice, Majority, and Right Shift operations

*/

module Miner(
	input clk,
	output out);
	//reg clk;
	reg done;
	reg [31:0] count;
	reg [639:0] header1, header2;
	reg [255:0] hashValues = 256'b0110101000001001111001100110011110111011011001111010111010000101001111000110111011110011011100101010010101001111111101010011101001010001000011100101001001111111100110110000010101101000100011000001111110000011110110011010101101011011111000001100110100011001;
	reg [2047:0] constantValues = 2048'b01000010100010100010111110011000011100010011011101000100100100011011010111000000111110111100111111101001101101011101101110100101001110010101011011000010010110110101100111110001000100011111000110010010001111111000001010100100101010110001110001011110110101011101100000000111101010101001100000010010100000110101101100000001001001000011000110000101101111100101010100001100011111011100001101110010101111100101110101110100100000001101111010110001111111101001101111011100000001101010011111000001100110111111000101110100111001001001101101101001110000011110111110111110010001111000011000001111110000011001110111000110001001000000110010100001110011000010110111101001001011000110111101001010011101001000010010101010010111001011000010101001110111000111011011111001100010001101101010011000001111100101000101010010101010000011000111000110011011011011000000000011001001111100100010111111010110010111111111000111110001101110000000001011111100111101010110100111100100010100011100000110110010100110001101010001000101000010100100101001011001110010011110110111000010101000010100101110000110110010000100111000010011010010110001101101111111000101001100111000000011010001001101100101000010100111001101010100011101100110101000001010101110111000000111000010110010010010111010010010011100100010110010000101101000101011111111101000101000011010100000011010011001100100101111000010010010111000101101110000110001110110110001010001101000111101000110010010111010000001100111010110100110010000011000100100111101000000111000110101100001010001000001101010101000000111000000011001101001001100000100010110000111100011011101101100000010000010011101001000011101110100110000110100101100001011110010110101001110010001110000001100101100110100111011011000101010100100101001011011100111001100101001001111011010000010111001101111111100110111010010001111100000101110111001111000101001010110001101101111100001001100100001111000000101001000110011000111000000100000100010010000101111101111111111111010101001000101000001101100111010111011111011111001101000111111011111000110011100010111100011110010;
	assign out = done;
	initial begin
	   count = 0;
	   done = 0;
	   header1 = 640'h0100000050120119172a610421a6c3011dd330d9df07b63616c2cc1f1cd00200000000006657a9252aacd5c0b2940996ecff952228c3067cc38d4885efb5a4ac4247e9f337221b4d4c86041b00000000;
	   header2 = header1; 
	   /*
	   clk = 0;
	   forever #10 clk=!clk;
	   */
	end
	Hash instance1(header1, hashValues, constantValues, status1);
	Hash instance2(header2, hashValues, constantValues, status2);
	always @ (posedge clk) begin
		if(count == 10000) done = 1;
		if(status1==1 & done==0) begin
		  count = count + 1;
		  header1[31:0] = {count[7:0],  count[15:8],  count[23:16],  count[31:24]};
		end
		else if(status2==1 & done==0) begin
		  count = count + 1;
		  header2[31:0] = {count[7:0],  count[15:8],  count[23:16],  count[31:24]};
		  end
		else done = 1;
	end
endmodule
